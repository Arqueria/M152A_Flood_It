module displayVGA(
    input wire CLOCK, //25 MHz
    input wire [2:0] BOARD [25:0][25:0],
    input wire [4:0] SIZE,
    input wire INITIALIZED,
    output reg [3:0] vgaRed,
    output reg [3:0] vgaBlue,
    output reg [3:0] vgaGreen,
    output reg Hsync,
    output reg Vsync
    
);



    


endmodule